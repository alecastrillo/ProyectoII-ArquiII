module adder (input logic [15:0] A,B,
										  output logic [15:0] out);
	assign out = A + B;	
	
endmodule 
