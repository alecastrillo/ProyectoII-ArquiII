module cmp (input logic [15:0] 	a, b,
				output logic 			out);
	
   assign out = (a==b);
	
endmodule 